module TOP(CLK, RST, IN);
  input CLK, RST, IN;

  SUB ccc(CLK,RST,IN);

endmodule

module SUB(input wire CLK,input wire RST,input IN, output OUT);
endmodule

