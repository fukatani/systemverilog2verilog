module TOP(CLK, RST, IN);
  input CLK, RST, IN;

  SUB ccc(CLK,RST,IN);

endmodule

module SUB(input  logic CLK,input logic  RST,input IN, output OUT);
endmodule

